library IEEE;
use IEEE.numeric_bit.all;

ENTITY testbench IS
END testbench;